LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY errorGenerator IS
PORT (
     );
END errorGenerator;

ARCHITECTURE makeError OF errorGenerator IS

BEGIN

END makeError; 
